* hongzhilian - 2FlipSynchronizer
.options post=2 list
*
* simulation time
.tran 1p 40n
*
* print list: clk, vin, Qm, Q
.print tran v(6) v(1) v(10) v(18)
*
.PARAM Vrail = 1.5V
.PARAM Tdelay = 13.1n
.PARAM TrL = 11.8n
.PARAM TrR = 13.8n
.global VCC
VCC VCC 0 DC Vrail
Vclk 6 0 PULSE(0 Vrail Tdelay 1n 1n 5n 10n)
Vin 1 0 PWL(0 0 TrL 0 TrR Vrail 14n Vrail 16n 0)
*
* instance inverters
XINV1 1 2 INV
XINV2 3 4 INV
XINV3 4 5 INV
XINV4 6 7 INV
XINV5 4 8 INV
XINV6 9 10 INV
XINV7 10 11 INV
XINV8 10 12 INV
XINV9 13 14 INV
XINV10 14 15 INV
XINV11 14 16 INV
XINV12 17 18 INV
XINV13 18 19 INV
*
* instance transmission gates
XTG1 2 6 3 7 TG
XTG2 5 7 3 6 TG
XTG3 8 7 9 6 TG
XTG4 11 6 9 7 TG
XTG5 12 6 13 7 TG
XTG6 15 7 13 6 TG
XTG7 16 7 17 6 TG
XTG8 19 6 17 7 TG
*
* define inverter
.SUBCKT INV IN OUT
M1 OUT IN VCC VCC mp L=1u W=20u
M2 OUT IN 0   0 mn L=1u W=20u
CL OUT 0.75p
.ENDS
*
* define transmission gate
.SUBCKT TG 1 2 3 4
M1 1 2 3 VCC mp L=1u W=20u
M2 1 4 3 0 mn L=1u W=20u
.ENDS
*
* details of the MOSFET model
.MODEL MP PMOS (level=2 LD=0.250U TOX=365E-10
+ NSUB=6.193910E+15 VTO=-0.826989 KP=2.2870E-05
+ GAMMA=0.4793 PHI=0.6 U0=241.796 UEXP=0.214214
+ UCRIT=19100.4 DELTA=0.859687 VMAX=47972.9 XJ=0.250U
+ LAMBDA=5.403347E-02 NFS=2.351269E+11 NEFF=1.001
+ NSS=1.0E+12 TPG=-1.0 RSH=76.020 CGDO=3.54775E-10
+ CGSO=3.54775E-10 CGBO=6.981174E-10 CJ=2.2624E-04
+ MJ=0.46650 CJSW=2.3825E-10 MJSW=0.24660 PB=0.700)
.MODEL MN NMOS (LEVEL=2 LD=0.250U TOX=365E-10
+ NSUB=2.13818E+16 VTO=0.84898 KP=5.7790E-05
+ GAMMA=0.8905 PHI=0.6 U0=610.8 UEXP=0.244555
+ UCRIT=128615 DELTA=2.0298 VMAX=92227.9 XJ=0.250U
+ LAMBDA=1.956049E-02 NFS=2.307838E+12 NEFF=1
+ NSS=1.0E+12 TPG=1.0 RSH=22.730 CGDO=3.54775E-10
+ CGSO=3.54775E-10 CGBO=6.354506E-10 CJ=3.7740E-04
+ MJ=0.45890 CJSW=5.1360E-10 MJSW=0.36620 PB=0.800)
*
.END